module main

import generator

fn main() {
	generator.create()
}
